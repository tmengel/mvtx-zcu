-------------------------------------------------------------------------------
-- Title      : mrDisc
-- Project    : ITS Readout Electronic Firmware
-------------------------------------------------------------------------------
-- File       : mrDisc.vhd
-- Author     : Piero Giubilato (piero.giubilato@cern.ch)
-- Company    : CERN
-- Created    : 2016-01-29
-- Last update: 2016-08-19
-- Platform   : Windows 10 64bit, Xilinx Vivado 2015.3
-- Target     : Xilinx Kintex-7 (XC7K325TFFG900-1)
-- Standard   : VHDL'2008
-------------------------------------------------------------------------------
-- Description: 'mrDisc' checks whether the 'INPUT' port had any rising edge
-- between two 'CYCLE' events (supposed to be in synch with 'CLK'), and outputs
-- a single '1' on 'OUTPUT' in synch with the 'CYCLE' signal and lasting one 
-- clock cycle if at least one rising edge has been detected, or a '0' otherwise. 

-- GENERICS: 
--   -> 'C_MRL' defines the level of Modulare Redundancy of the hardened components
--      should be odd and it is anyway suggested to only use the 3 and 5 values. 
--      The 'INPUT' port width is equal to 'C_MRL'. 
--   -> 'C_MRO' defines wheter the modular redundancy stops at the port output
--      ('C_MRO = false'), in which case the output is a single bit port, or when
--      the modular redundancy is carried outside the entity ('C_MRO = true'), in
--      which case the 'DIFF' port is a parallel bus 'C_MRL' wide of fully
--      triplicated circuits. The 'OUTPUT' port width is equal to 'C_MO'.
--
-- I/O PORTS:
--  ->  'CLK' is the entity clock, and the outputs are synchronous with this clock,
--      i.e. they change state just after the 'CLK' rising edge.
--  ->  'RST' is the active-high synchronous reset. The unit start working after
--      'RST' goes low.
--  ->  'EN' active high enable, if low forces the output to '0' (no transition
--      signalled whichever the input). This input is asynchronous.
--  ->  'CYCLE' is the input for the pattern cycle, should be in synch with the clock,
--      and asserted at every pattern cycle end.
--  ->  'READY' is the input for the pattern status, should be in synch with the 
--      clock, and asserted at every pattern cycle end. Transition on the 'INPUT'
--      signal are recorded only when 'READY = 1'.
--  ->  'INPUT' is input signa, 'C_MR' replicated.
--  ->  'OUTPUT' is the output, asserted in synch with 'CYCLE' and equal to '1'
--      in case a rising edge has been detected during the interval between the last
--      and the current 'CYCLE, '0' otherwise. The '1' level remains asserted for 
--      one clock cycle only.
--  ->  'WARN' is a warning flag which if '1' indicates that within the comparator
--      voting system not all signals agree, i.e. that some upset is affecting the
--      comparator itself. The signal is synchronous with 'CLK' and tied to '0' 
--      during reset.
--

-- Libraries.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- Packages.
use work.mrTools_pkg.all;


--------------------------------------------------------------------------------
--                             Entity Declaration                             --
--------------------------------------------------------------------------------
entity mrDisc is
    generic (
        C_MRL:   natural := 3;       -- Modular Redundancy Level.
        C_MRO:   boolean := false    -- Modular Redundancy Output.   
    );
    port (  
        CLK:    in  std_logic;
        RST:    in  std_logic;
        EN:     in  std_logic;
        CYCLE:  in  std_logic;
        READY:  in  std_logic;
        INPUT:  in  std_logic_vector(C_MRL - 1 downto 0);
        OUTPUT: out std_logic_vector(mrPortWidth(1, C_MRL, C_MRO) - 1 downto 0);
        WARN:   out std_logic
    );
    
    -- Make 'rtDisc' untouchable by the synthesis/placement tools. 
    attribute DONT_TOUCH of mrDisc: entity is "TRUE";
        
end mrDisc;

--------------------------------------------------------------------------------
--                     Architecture 'Behavioral' Declaration                  --
--------------------------------------------------------------------------------
architecture Behavioral of mrDisc is

    -- Output signals generated by C_MRL replicated discriminators.
    signal sDsc: std_logic_vector(C_MRL - 1 downto 0):= (others => '0');    
        
begin
    
    -- Discriminators, 'C_MRL' replicated. Compares the 'SIG1' and 'SIG2' inputs
    -- and asserts a '1' if they differ. Purely async process.
    MR: for i in 0 to (C_MRL - 1) generate
        DSC : entity work.muDisc
        port map (
            CLK    => CLK,
            RST    => RST,
            EN     => EN,
            CYCLE  => CYCLE,
            READY  => READY,
            INPUT  => INPUT(i),
            OUTPUT => sDsc(i)
        );
    end generate MR;
        
    -- Output voting stage. Votes the values of the 'C_MRL' 'rDiff' registers,
    -- and directly drives the 'OUTPUT' and 'WARN' ports.
    MR_VOTE: entity work.mrVotingStage
    generic map (
        C_WIDTH => 1,
        C_MRL => C_MRL,
        C_MRO => C_MRO
    )
    port map (
        INPUT   => sDsc,
        OUTPUT  => OUTPUT,
        WARN    => WARN
    );
    
end Behavioral;
