-------------------------------------------------------------------------------
-- Title      : watchdog
-- Project    : RUv1
-------------------------------------------------------------------------------
-- File       : watchdog.vhd
-- Author     : Arild Velure <arild.velure@cern.ch>
-- Company    : CERN European Organization for Nuclear Research
-- Created    : 2016-04-28
-- Last update: 2017-09-27
-- Platform   : Xilinx Vivado 2017.4
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: wishbone watchdog
-------------------------------------------------------------------------------
-- Copyright (c) 2016 CERN European Organization for Nuclear Research
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2017-02-07  1.2      AV      Converted from watchdog.sv
-------------------------------------------------------------------------------
--
-- Currently can not be used as the RUv1_testbench.sv forces the input timeout_i input 
-- from the testbench, but Cadence does not support forcing VHDL signals from SV, so 
-- this module must be written in SV. Use watchdog.sv instead.
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity watchdog is
  generic(
    TIMEOUT_BIT_WIDTH : natural := 16
  );
  port(
    clk_i          : in  std_logic;     -- clock input
    rst_i          : in  std_logic;     -- synchronous reset input

    stb_i          : in  std_logic;     -- strobe input
    cyc_i          : in  std_logic;     -- cycle input
    err_o          : out std_logic;     -- error output

    actual_state_i : in  std_logic_vector(TIMEOUT_BIT_WIDTH - 1 downto 0); -- 
    actual_state_o : out std_logic_vector(TIMEOUT_BIT_WIDTH - 1 downto 0); -- 
    timeout_i      : in  std_logic_vector(TIMEOUT_BIT_WIDTH - 1 downto 0) -- timeout value
  );
end entity watchdog;

architecture RTL of watchdog is

  signal s_transaction_active : std_logic;
  signal s_counter            : std_logic_vector(TIMEOUT_BIT_WIDTH - 1 downto 0);
  signal s_rst_cntr           : std_logic; -- resets the upcounter
  signal s_is_equal           : std_logic;

begin
  s_transaction_active <= cyc_i and stb_i;

  INST_timeout_upcounter : entity work.upcounter_core
    generic map(
      BIT_WIDTH     => TIMEOUT_BIT_WIDTH,
      IS_SATURATING => 0,
      VERBOSE       => 0 )
    port map(
      CLK            => clk_i,
      RST            => rst_i,
      RST_CNT        => s_rst_cntr,
      CNT_UP         => s_transaction_active,
      CNT_VALUE      => s_counter,
      ACTUAL_STATE_O => actual_state_o,
      ACTUAL_STATE_I => actual_state_i);

  s_is_equal <= '1' when (s_counter = timeout_i) else '0';
  s_rst_cntr <= '1' when (s_transaction_active = '0') else s_is_equal;
  err_o      <= '0' when (s_transaction_active = '0') else s_is_equal;

  -- synthesis translate_off
  p_assert_timout : process(clk_i) is
  begin
    if rising_edge(clk_i) then
      assert (err_o = '0') report "Timeout generated by wishbone Watchdog!" severity WARNING;
    end if;
  end process;
  -- synthesis translate_on
end architecture RTL;
